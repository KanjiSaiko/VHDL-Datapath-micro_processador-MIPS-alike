library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity processador_MIPS is
	port (
		clock	: in std_logic;
		reset	: in std_logic
        --Reg_out    : out std_logic_vector(7 downto 0)
		);
end processador_MIPS;

architecture behavior of processador_MIPS is

    signal PC	: std_logic_vector(7 downto 0); -- Contador de programa (Program Counter) que armazena o endereço atual de execução.
    type mem_dados is array (integer range 0 to 255) of std_logic_vector(7 downto 0);
    type mem_instruc is array (integer range 0 to 255) of std_logic_vector(15 downto 0);
    type banco_regs is array (integer range 0 to 15) of std_logic_vector(7 downto 0);

    signal mem_i    	        : mem_instruc:= ( --Memória de Instruções, com 255 posições de 16 bits cada.
        0 => "0000000000000001", -- LDA endereço 1 para R0
        1 => "0000000100000010", -- LDA endereço 2 para R1
        2 => "0011001000000001", -- ADD R0 + R1 -> R2 => 4
        3 => "0111001000000001", -- STA R2 no endereço 1
        others => (others => '0') -- Demais posições zeradas
    );

    signal mem_d	            : mem_dados := ( --Memória de Dados, com 255 posições de 8 bits cada.
        0 => "00000000",
        1 => "00000001", --1
        2 => "00000011", --3
        others => (others => '0') -- Demais posições zeradas
    ); 

    signal regs                 : banco_regs := (others => (others => '0')); --Banco com 16 Registradores
    signal desvio	            : std_logic; --Controle para indicar se deve ocorrer um salto (branch).
    signal opcode  	            : std_logic_vector(3 downto 0); --Código de operação das instruções.
    signal ula		            : std_logic_vector(15 downto 0); --Saída da ULA que executa operações aritméticas.
    signal equal	            : std_logic; --Sinal para verificar se R0 é igual a R1 (usado em instruções de comparação).
    signal instrucao	        : std_logic_vector(15 downto 0); --PEGA A INSTRUÇÃO DA POSIÇÃO ATUAL
    signal enable_reg	        : std_logic; --Habilita a gravação de valores em registradores.
    signal R0, R1               : std_logic_vector(7 downto 0);

begin --a memória de instruções é carregada com valores iniciais. Cada posição contém uma instrução.
    
    

    enable_reg	<= '1' when (opcode = "0000") or (opcode = "0001") or (opcode = "0010") or (opcode = "0011") else
				'0';

    --Verifica se R0 e R1 têm valores iguais.
    equal <= '1' when (R0 = R1) else
        '0';

    --Indica se um salto deve ocorrer.
    desvio <= '1' when (opcode = "0100" and equal = '1') or (opcode = "0101" and equal = '0') or (opcode = "0110") else
        '0';

    

    process(reset, clock)
        begin
            if (reset = '1') then   --Se reset está ativo (1), ele zera tudo
                R0	 <= (others => '0');
                R1   <= (others => '0');
                regs <= (others => (others => '0'));
                PC   <= (others => '0');

            elsif (clock = '1' and clock'event) then
                -- LEITURA DA INSTRUÇÃO
                instrucao <= mem_i(conv_integer(PC));
                opcode <= instrucao(15 downto 12);

                if(enable_reg = '1') then
                    R0 <= regs(conv_integer(instrucao(7 downto 4)));
                    R1 <= regs(conv_integer(instrucao(11 downto 8)));
                end if;

                -- Decodificação e execução
                case opcode is
                    when "0000" => -- LOAD
                        regs(conv_integer(instrucao(11 downto 8))) <= mem_d(conv_integer(instrucao(7 downto 0)));
                    
                    when "0111" => -- STORE
                        mem_d(conv_integer(instrucao(7 downto 0))) <= regs(conv_integer(instrucao(11 downto 8)));
                    
                    when "0001" => -- ADD
                        ula <= regs(conv_integer(instrucao(7 downto 4))) + regs(conv_integer(instrucao(11 downto 8)));
                        regs(conv_integer(instrucao(11 downto 8))) <= ula;

                    when "0010" => -- SUB
                        ula <= regs(conv_integer(instrucao(7 downto 4))) - regs(conv_integer(instrucao(11 downto 8)));
                        regs(conv_integer(instrucao(11 downto 8))) <= ula;

                    when "0011" => -- MULT
                        ula <= regs(conv_integer(instrucao(7 downto 4))) * regs(conv_integer(instrucao(11 downto 8)));
                        regs(conv_integer(instrucao(11 downto 8))) <= ula(7 downto 0);

                    when others =>
                        ula <= (others => '0'); -- Valor padrão

                    end case;

                if (desvio = '0') then --Se não houver desvio.
                    PC <= PC + 1;

                else --Caso contrário, ele pula para o endereço indicado. --JUMP, BEQ OU BQE
                    PC <= PC + instrucao(7 downto 0);
                end if;
            end if;
                    
            end process;
end behavior;